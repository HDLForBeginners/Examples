`define VERSION_MAJOR 1
`define VERSION_MINOR 1
